// includes everything
// cores
// llc
